module test;
  initial begin
    $display("Hello, simulation!");
    $finish;
  end
endmodule
